`ifndef __RSA_DEFINE__
`define __RSA_DEFINE__

parameter RSA_MAX = 1024;
parameter RSA_BUS = (RSA_MAX-1);
parameter RSA_MAX_LOG2 = 12;

`endif